--------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:	00:43:56 09/28/2013
-- Design Name:
-- Module Name:	C:/Users/fadeev/Documents/dmkonsttdt4255_work/hardware/sign_extender_tb.vhd
-- Project Name:	exercise1_mux_work
-- Target Device:
-- Tool versions:
-- Description:
--
-- VHDL Test Bench Created by ISE for module: sign_extender
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes:
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.	Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;

ENTITY sign_extender_tb IS
END sign_extender_tb;

ARCHITECTURE behavior OF sign_extender_tb IS

		-- Component Declaration for the Unit Under Test (UUT)

		COMPONENT sign_extender
		PORT(
				input : IN	std_logic_vector(15 downto 0);
				output : OUT	std_logic_vector(31 downto 0)
				);
		END COMPONENT;


	--Inputs
	signal input : std_logic_vector(15 downto 0) := (others => '0');

	--Outputs
	signal output : std_logic_vector(31 downto 0);
	-- No clocks detected in port list. Replace <clock> below with
	-- appropriate port name

	constant clk_period : time := 10 ns;

BEGIN

	-- Instantiate the Unit Under Test (UUT)
	uut: sign_extender PORT MAP (
					input => input,
					output => output
				);

	-- Stimulus process
	stim_proc: process
	begin
			-- hold reset state for 100 ns.
			wait for 100 ns;
			-- insert stimulus here

			wait for clk_period*10;
			input <= ( others => '0');

			wait for clk_period*10;
			input <= ( others => '1');

			wait for clk_period*10;
			input <= "0101101110100010";

			wait for clk_period*10;
			input <= "1111010001011011";

			wait;
	end process;

END;
