-- blablabla