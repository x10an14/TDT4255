----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:	15:01:07 09/20/2013
-- Design Name:
-- Module Name:	simple_multiplexer - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity simple_multiplexer is
generic (N :NATURAL);
	Port(
		a : in  STD_LOGIC_VECTOR (N-1 downto 0);
		b : in  STD_LOGIC_VECTOR (N-1 downto 0);
		control_signal : in  STD_LOGIC;
		output : out  STD_LOGIC_VECTOR (N-1 downto 0));
end simple_multiplexer;

architecture Behavioral of simple_multiplexer is

begin
	output <= b when control_signal = '1' else
				a;

end Behavioral;
